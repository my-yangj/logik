//env.sv
